<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-18.4917,0.256351,103.908,-60.2436</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>6.5,-8.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>6.5,-16.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>25,-12</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>29,-12</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>7.5,-11.5</position>
<gparam>LABEL_TEXT AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>CC_PULSE</type>
<position>-40.5,-11.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>6.5,-24.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>6.5,-31.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>21.5,-27.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>25.5,-27.5</position>
<input>
<ID>N_in2</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>7,-28</position>
<gparam>LABEL_TEXT OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>6.5,-47.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>6.5,-39.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AO_XNOR4</type>
<position>-70.5,-37.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>30</ID>
<type>BA_NAND4</type>
<position>22.5,-43.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>32</ID>
<type>AO_XNOR4</type>
<position>-35,-35</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>27,-43.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND4</type>
<position>-45,-48.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>5,-42</position>
<gparam>LABEL_TEXT NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>76.5,-12</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AO_XNOR2</type>
<position>76.5,-27</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>BE_NOR2</type>
<position>78,-44</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>55.5,-9.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>48</ID>
<type>CC_PULSE</type>
<position>26.5,-1.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>55.5,-15.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>51,-25</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>51,-32</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>51,-40.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>51,-49</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>80.5,-12</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>80.5,-27</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>82,-44</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>49.5,-12</position>
<gparam>LABEL_TEXT xorgate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>49,-27.5</position>
<gparam>LABEL_TEXT x nor gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>49.5,-43.5</position>
<gparam>LABEL_TEXT nor gaTE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-11,15,-8.5</points>
<intersection>-11 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-8.5,15,-8.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-11,22,-11</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-16.5,15,-13</points>
<intersection>-16.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-16.5,15,-16.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-13,22,-13</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-12,28,-12</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>8.5,-24.5,18.5,-24.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>18.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>18.5,-26.5,18.5,-24.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-24.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-31.5,13.5,-28.5</points>
<intersection>-31.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-31.5,13.5,-31.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-28.5,18.5,-28.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-28.5,25.5,-27.5</points>
<connection>
<GID>20</GID>
<name>N_in2</name></connection>
<intersection>-27.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-27.5,25.5,-27.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-40.5,13.5,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-39.5,13.5,-39.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-40.5,19.5,-40.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection>
<intersection>16.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-42.5,16.5,-40.5</points>
<intersection>-42.5 6</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16.5,-42.5,19.5,-42.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>16.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-47.5,13.5,-44.5</points>
<intersection>-47.5 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-47.5,13.5,-47.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-44.5,19.5,-44.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>13.5 0</intersection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-46.5,19,-44.5</points>
<intersection>-46.5 4</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-46.5,19.5,-46.5</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>25.5,-43.5,26,-43.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-43,64,-40.5</points>
<intersection>-43 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-43,75,-43</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-40.5,64,-40.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-49,64,-45</points>
<intersection>-49 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-49,64,-49</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-45,75,-45</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-32,63,-28</points>
<intersection>-32 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-28,73.5,-28</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-32,63,-32</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-26,63,-25</points>
<intersection>-26 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-25,63,-25</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-26,73.5,-26</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-11,65.5,-9.5</points>
<intersection>-11 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-11,73.5,-11</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-9.5,65.5,-9.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-15.5,65.5,-13</points>
<intersection>-15.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-15.5,65.5,-15.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-13,73.5,-13</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-27,79.5,-27</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-44,81,-44</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>64</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>